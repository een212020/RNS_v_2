`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 05.04.2023 21:11:01
//////////////////////////////////////////////////////////////////////////////////


module FA(
    output Cout, Sum,
    input A, B, Cin
    );
    assign Sum = A^B^Cin;
    assign Cout = A&B | B&Cin | Cin&A;
endmodule
